��   �`]                                                                                                                                                  ��                                                                      �����                                                                      ����                                                                     ����                                                                    ����                                                                   ����                                                                   ���                                                                   ���                                                                  �����                                                        ����                                                     ����                                                   ����                                                ����                                               X�����                                              ����                                               ����                                               ����                                               �����                                              ������                       ѡ                        ����                         ѡ�                     ��������                           ��Y            �������                            �鉊AA   ������                             ����鈠YX�����������                              ���������҈�XYY����AAA����                              ���������щYZY���ꠈ���BBBA�����                               ���������ш�AXYX���ъ�+++A�������                               �������҈���AABXX�   ��*++*�����                               �������顡���AAAX���  ь*+****���                               ������҈������X@���  �++++**���                                ���������������@��s++++**��                                �AAA�������������AA�++++++*�                                AAAAAAAA�����������AA++++++++*���                                 �AABAABBYXA������������**++++++ss�                                  �@ABBBBBYY���҈������*+++++*ss�                                  �@AAAAABY����҉����+++++sr�                                   С��AAAABB���҉����***+++*s�                                     ������AAAA��Ӊ������***+++*s�                                       щ������AAAA��������**+*r                                       щ����AAAAAA�������***��                                          鉊��AAAAA��������**r                                             �ꉡ�AAA�������ss�                                               鉊�@�������ssssr                                                   ꉊ������������sssssr�                                                     鈉������҈�ssssssr                                                       �뉡�����sssssss�                                                           ��sssssss�                                                                 �ss�                                                                 s++**�                                                                 ++++**+*�                                                                ++++++++++�                                                                �++++++++++                                                                �*+++++++++                                                                 *+++++++                                                                 �+++++++                                                                  Ҋ*++++++�                                                                  �s*+++++�                                                                  s*+++++�                                                                  r*++A�                                                                   ъ���                                                                    ����                                                                    ���                                                                    ���                                                                     ���                                                                     ���                                                                     ꣤�                                                                     ��                                                                     ���                                                                     �����                                                                      ����                                                                      �舉��                                                                      鈉��                                                                     ������                                                                     ������                                                                     ������                                                                      뉊���                                                                      �����                                                                       щ���                                                                       늡�                                                                       艡�                                                                       ����                                                                        鉣                                                                        ��                                                                         顠                                                                         ��                                                                        ъ�                                                                        ���                                                                      ����                                                                     ����                                                                   ����                                                                                                                                        �                                            