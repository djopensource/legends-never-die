��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                                                            ��                                                            ��                                                            ����                                                       ꉉ�� ��                                                      뉉��� ꠠ���                                                      늡��  頉���                                                       ��������                                                         �AABBBX����                                                     ��AABBBBBBBX���                                                 ѡ�AABXXBBBBBBX���                                              �AABXYXAAABY@��                                             �AABXYX       χ��                                     �BBBBB       ��                                     ABBBA�      ���                                      AAA��    ���                                      A���  X���                                        AA������A��                                         �������                                          �@@��������                                            ꣤@@@���҉������                                              ��������҉������                                              ���������ш����                                                �������������щ���                                                 ���������������� Љ����                                                   �����������������                                                        ң��������������                                                          �������������҈�                                                           ���������������                                                            늋������������                                                            ��������������                                                             ���������                                                             ����                                                            ����                                                            ����                                                            ���++***r                                                          �++++++++++++**�                                                          �++++++++++++Ћ+�                                                        �++++++++++++*rӌ+�                                                       �+++++++++++**Ҋ*++s                                                      �+++++++++++++*sщ*++s                                                     +++++++++++++++҉*++s                                                    +++**+++++++++++�ӌ+*s                                                   **********++++�ӌ+�                                                  �������*++++�Ҍ*�                                                 sssss����ssss�*+***��*                                                �ssss�������sss*****��*�                                                �sr��� �s�***s��                                               ssr���   싋ts��                                              sssr��     �s�ь��                                              �ssss��       �������                                             �ssssr�        ӊs������                                            ��sss���           Ԋ����������                                            �������             ꉊ�������                                           �������               舉�������                                           ������                 鉊������                                        �����                    ������                                       Z����                   �AAA��                                      YYBA����                   BBAA��                                      YBAA��                    XBBA��                                      YYBBA��                    YBBA�                                     �YXBA��                     XYBA��                                     YBBA�                      BBBA���                                     BBBAA�                       BBA��                                    BAA��                      AA���                                     �YBA��                       AAA���                                    BA��                        AAA��                                    BAA��                         AA���                                     BA�                          AA��                                    �BA�                          AA���                                    A��                           A��                                    �A�                            A��                                    ����                             ��                                   ��                             A�                                   ��                            A��                                   �����                           A��                                   �������                          ��                                   ꉉ���鉢��                     ����                                                               �������                                                                 ������                                                            렡�������                                                               �������                                                                                                                                                              