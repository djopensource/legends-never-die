��   �2�l                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �����                                                                                                     ��                                                                                                   ����                                                                                                   ���                                                                                                  ꡤ����                                                                                                  ꉊ������                                                                                                 �ꉊ������                                                                                                 Ѣ��                                                                                                  졡�����                                                                                                 ����������Ѣ                                                                                                 ������                                                                                                  ѡ��Ѥ                                                                                                  ѡ���ң                                                                                                  ������                                                                                                   ����                                                                                                    ��������                                                                                                     ��������                                                                                                      ��������                                                                                                       ꡊ���                                                                                                        ������                                                                                                        Ҋ���                                                                                                         Ҋ�                                                                                                         �щ�����                                                                                                         鉉�ԡ���                                                                                                         룤��                                                                                                        ꊣ���                                                                                                        ъ�����                                                                                                        ъ��                                                                                     �          ъ��       ꡣ�                                                                      �����       ��ѡ��   ���                                                                 �������  顢�������������������                                                            ��������������������������������������                                                         颢��������������������������������������                                                      ����������������������������������������                                                    �����������������������                                                 �������������������XAAA                                               ��BX���������������X�                                           �AA��������A����                                       �������������������                                    ���Ҋ��������������                                 ��������B����������                              顤��Ҋ��������������                          ꢤXX���Ҋ��A���������������                       ��AXX�������A���������������                      좤A��������������҈�����ӈ��Ң                    ꡤAAXXX��Y����XX�   ���҈������ꈉ���                  ꡢ�XX��������        �ꉊ������ꈈ����                顋�������X�            艉��������҈��              ꡢ������   �A���              ������ӈӈ���            衡��������     ��                   ���ӈӈ����          �������A����        �A�                     �����ӈ����          ���������           �����                       ����ӈ���        ����������              ��X��                         ����뉊���        ����������                 ҢX���XX                         ��҉�����        ����������                 �X���X                          �鈉���        ���������                  �Y���X                           �鉢        ��������                  �X����XXXX�                            �鉣       ��������                    �X�����X�                             ��       ������                    �������XXZX�                            ��      �������                      �Ҋ�����XXXYY�                                  ������                      ��щ����XX�                           �X     ������                       ��҉����XX                           щXA      �����                    �щ�����                            XAAA      늊�������                   �ꊣ�                             �XA       ���������                  �ш��                             XX�        ������������                 ��뉢�                              �X         �������������                 鉉�                               ��X�         뢊�����������                  �ꉡ                                �          ������������                  �҉���                                  �            �����������                   ҉��                                    ��             銉���������                    �늤��                                                     ���ӈ����                    �슣�                                                         ���������                      뉡����������������������                                                                                                                                                                                                                                                                                                                                                                                                                �   ����   ���  ���   ��   ���   ���       ��  ���  ��  ���   ����       ��   �� ���         �   �  �� ��  �ꤢ  ��  �        ��  �   ��� ��  ���       롡�  � ��         �   �    �  ��   �� ��  �         ��      �� �    ���       �  � ��          �   �    �    ��   �� ��  �         ��      � �    ���       �  � ��          �   �    � ��   �� ��  �         ��  �     � �   ���       �  � ��          �   ��  ��� ��  �� ��  ���       ��  ��   ��  ��  ��        �  � ���         �   �  �� ��  �� ��  �       ��  �    �  �  ��       �  � ��         �   �    �� ��   �� ��    �       ��       ��  �    ���       �  � ��          �   �    �� ��   �� ��     �       ��       ��  �    ���       �  � ��          �   �    �� ��   �� ��     �       ��       �  �    ���       �  � ��          �  �  �� ��  �� ���  ���       ��  �    �  ��  ���       롡�  � ��         뢢�  ����  ����  ���   ���   ��   ���       ���  ���       ���   ���       ��   ��  ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            