��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         �                                                                                                                                                                                                       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      衢�                                         ��                                      ����                                       ���                                       ���                                       ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �                                                                                                                      �                                                             X�                                                             XW                                                             �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          