��   |pd                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��                                                         Ј��                                                        Ҋ����                                                     �����oo                                                   �������                                                ������                                 �������  ��������                                ��������������щ��XB��������                                 YXAA����������������ш�XYYXBA��������                                 ZXAA����������������҈�ABAAA������                                  YYBAAA����������������҉�AA������                                     AAAAA@�������������Ј�������                                        AAAAAA������������ш��������                                          A@A@@�������������щ����                                             �@�����������ꈈ�����                                                 �������������銊����                                                 �������ӈ��������                                                  ��������ӈ���ꢢ��                                                   �������ш����룢�                                                  ����щ���衡���                                                   �����щ�����늢���                                                   �����������o�Љ������                                                    ��������q���������                                                    �������ꈈ�������                                                    ���������������������                                                     �������������҈����҈���                                                     ъ����������������������                                                     Ҋ����������������������                                                      ъ��������҉�����������                                                      ���������҉�����������                                                        �� ����ш����������                                                            �����ш����������                                                            ��ш�������������                                                            ��ш�������������                                                           ъѺш��҉���������                                                          ��Ѻш��҈��������                                                          �rqш������������                                                          �ssr������������                                                         �����������                                                         �**�                                                          �*+++**�                                                          �s*+++++**�                                                          �s+++++++++*�                                                           ��s*++++++++*                                                           ��s**+++++++*�                                                            ��r**++++++++�                                                             ���*++++++++�                                                              ����s*+++++++A�                                                               Ӻ�s*+++++BB                                                               ����*++AABX                                                                �r���s*@AAAA                                                               �rr���s��AAAA�                                                              ���rr�ъ��AAAA                                                             ���rrsӉ����AAA                                                            ���rrrӈ�����@AX                                                            л�rssr������A                                                           �ѻ�ssss���������                                                          ��кrss�щ������                                                         ����r���  �������                                                          ����҉�   Њ�����                                                         �����҉�   ������                                                     �����҉   Ѣ�����                                                   �XAA�����҈   ����                                                   �AAA��������   ���                                                 ����������   ���                                               ��������������    ���                                              ����������     �������                                           ���������            �������                                         �����������               늣����                                       ��������                  Ҋ�����                                       �����                     ������                                      ������                        늋���                                       颤����                          ъ����                                      ꠢ���                          �����                                        ����                          늊��                                         ���                         Ҋ���                                          ����                        щ���                                           頣�                       ����                                           ���                      �����                                            щ�                        ꉊ��                                                                         Љ���                                                                        뉊��                                                                        �Ӊ��                                                                       ��뉉�                                                                     �������                                                                   �������                                                                  ������                                                                   �����                                                                                                                                                                                        