��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                                                             ꉠ��                                                              Ј����                                                             ���������                                                             ���������                                                            ���������                                                              Љ����ꉉ���                                                              ����ш����                                                              ���ш���                                                              Љ�AAX                                                                �AAXYYXXY�                                                              �AAXYZZZYYY�                                                            �XABXYYZZZYYYY�                                                          XAAABXYYZZYYXX                                                         BAAAAAAAABBBBAAA�                                                 � BAAAAA@@AAAAAAAA�                                                 ����AAAA@@@@@AAAAAAA�                                                ѡ��AAA@@@��AAA@AA�                                                ����AAAAAA@����@@��                                                �뉉�@AAAA@�������@@�                                                �щ��뉤@AAAA@��������                                                   ��Ј�AAAAAAA����������                                                      Ј�AAAAAA����������                                                       ЉAAAAAA���������                                                         СAAAAAA���������                                                          �AAAAA���������                                                           ФAAAA@���������                                                          �AAAA@���������                                                        AA��@���������                                                      �AA@������������                                                     AA���������������                                             BA�����������������                                        Ј��A������������������                                        ���������룤������AA�                                      ��������Ѣ������@@�����                                      ����       Њ�������**++�                                     ω����         ҋ*++++++++��                                               s*****++++++++++�                                                       s+*�*++++++++++�                                                      �*+�r++++++++++�                                                      ��++++�ԉ*+++++++++�                                                    �+++++��s**++++++**+�                                                   �+++++���r**+++++*�                                                 �+++++����t*******��                                                �+++*���s*++***sss�                                              Ԍ++*����******srrsss��                                             �++++*���s*****�srrrsrrs�                                            �++++��**�ssr�rssss�                                           �AB++���rsss�Ѻ�rrsss                                          AAAA���sts��  �ssss                                         AAA���ss�    �ssss                                        ���ts��      Ӌsss                                       ��������ss��        ҋ�ssss�                                      ����������          ��s�����                                      �������               ъ������                                      ������                 �������                                      ������                    뢡����                                      ꊣ�                     �������                                       ��A�                     ъ����                                       ꢤAA�                     ����AB�                                     ��AA�                      ��AAXX                                    ���AA                      �AABYY                                    ꣤AA�                       �ABBY�                                   ��A�                        �ABBBX                                  ���                         �ABBA�                                  ����                          ѤAAAAA�                                  ң��                           �A�                                  ���                           ꊣAA�                                 ���                             �AA�                                  룤�                              ңAA�                                 Т��                               �AA�                                 ���                                �AA�                                 ��                                ���                                 ѣ�                                ���                                Ѥ�                                 ���                               ѤA�                                  뢣                               �AA�                               颣�                             �AA                            ����                           ����                            ��������                         ��                                �����                      A�                                  ��                     ��                                                             �����                                                                ��                                                           