��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           鉢�                                                            Ҋ����                                                            �����                                                             ��뉡�                                                            艊�����                                                             ҉��������                                                             �����������                                                             ����҈���                                                           ������                                                         ZXYZYXB��                                                          �ZZZYXXY�                                                            YYYZZZZYXBY                                                          YBBYZZZYYYYBBY                                                         XBABBXBBAAAAABAXZ    �                                               �AAAAAAAAAAAAAAABY ѣ�                                               �AAAAAAAAAA@AAAAAAB���щ                                             �AAAAAA@��AAAAAAA���Ѣ                                              �@@���AAAAA����ѡ�                                             �@@�������AAAAAA������                                              �@��������AAAA@���                                                  �����������AAAAA����                                                    ������������AAAAA�                                                     ������������AAAAA�                                                        Ӌ����������@AAAA�                                                        Њ����������@AAAA�                                                        �����������@AAAA�                                                         ������������@AAAA�                                                          щ����������AAAY                                                         �����������@@ABX                                                      ���������������AAB�                                                   ���������������AA�                                            ������������������AAB��                                     �����������뉉�������                                    ӌ�������������� ��ꈉ������                                  A++*++++++*ss��      ���                                  +++++++++++*�           �ψ�                                   �+++++++++++*r��                                                 �++++++++++++*sҌ**s                                                       �+++++++++++++щA+++�                                                     �++*+++++++++++��ӌ+++s                                                    �+***++++++++++sыB�                                                  �***+++++++++���A+++�                                                 �ss*+++++++++�ь+++s                                                s��rrs�*++++++++sҋ++++s                                              rssss���ss�*++++++sы+++++�                                             �s��s������sss*++++*sъ+++�                                            sssssssrr����ss**++*sЉ*+++B�                                           �s��sssrs�   �s�***sЉ*BBB�                                           Ԋ�sssss��    �Ԋ�sӣAA�                                          �ssssss��       Ԋ���                                         ҉ssssss��         Ԋ������������                                        �ԉ�����           ҉����������                                        �����뉉             ꉡ�������                                       �����                  늉����                                       ���뉠                    ������                                     ����                    A���                                      ����                    �AA����                                      XA���                    �AA���                                      YA��                     AA���                                     XBA��                     �AAA���                                      BAA�                     �A���                                      �AAA�                    ������                                      A�                     ����                                      A���                      ����                                       AA��                       ����                                      A�                        ����                                       A��                         �����                                       ���                         ���                                       A��                         ��                                       �                         ��                                       ��                          ��                                       ���                          ���                                      ��                         ��                                      ���                          ��                                       ��                       ��                                     A��                     �����                                      ������                   ����                                                               ����                                                                    �����                                                                      �                                                                     �                                                                      �                                                                                                                                                                     