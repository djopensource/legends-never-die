��   �`]                                                                           ��                                                                       衡��                                                                      顡�                                                                      щ��                                                                     鉣�                                                                     щ��                                                                      ꉢ                                                                      ꉡ                                                                     ꉠ��                                                                    �ꉢ                                                           舠��                                                        �ꉢ                                                     �ꈠ                                                  �ꈊ�X                                                  ꉡ�                                                 鉡�                                                 ꊣ�                                                 ꢣ��                                                 ꠣ����                                                 늢�                        ��                           좢�����                     ���                            �������            Y���                             ������   AA����                              ������戈���XY�������                               늢�AAA����YYX������������                                �����ABBB������銣YZY��������щ�                                Љ�����A+++������XYXA��������ш��                                 ꉉ��*++*��   �XXBAA���������ҡ�                                ꉉ****+*��  ꈈXAAA���������ш��                                ъ�**++++�  Ј�@X��������҈����                                ��**++++sԊ@���������������                                 �*++++++�AA�������������AAA�                                  ъ�*++++++++AA�����������AAAAAAAA                                  �ss++++++**������������AXYBBAABAA�                                  �ss*+++++*��������҉�YYBBBBBA@�                                   �rs+++++�������҈�YBAAAAA@��                                     �s*+++***�������ҊBBAAAA����                                      �s*+++***�������Ӊ�AAAA������                                      r*+**��������AAAA��������                                        ��***�������AAAAAA������                                         r**��������AAAAA�����                                           �ss�������AAA�����                                              rssss�������@����                                                �rsssss���������������                                                   rssssss���Ӣ�������                                                      �sssssss��Ӊ�����                                                        �sssssss��                                                           �ss�                                                                 �**++s                                                                 �*+**++++                                                                 �++++++++++                                                                ++++++++++�                                                                 +++++++++*�                                                                 +++++++*                                                                 +++++++�                                                                 �++++++*��                                                                  �+++++*s�                                                                  �+++++*s                                                                  �A++*r                                                                   �����                                                                    ����                                                                    ���                                                                    ���                                                                    ���                                                                     ���                                                                     ����                                                                     ���                                                                     ����                                                                     �����                                                                     ����                                                                      ꊉ���                                                                     �����                                                                     ꤡ���                                                                     ������                                                                     ������                                                                     ������                                                                      �����                                                                      �����                                                                      ����                                                                      ����                                                                       ꣊�                                                                       ���                                                                        ��                                                                        ���                                                                        ��                                                                        ���                                                                       ���                                                                       ����                                                                      ����                                                                     ����                                                                                                                                               �                            