��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ����                                                            ꉊ���                                                             Љ�����                                                            �������                                                            ��������                                                            颣�������                                                              �����������                                                              늊�҈���                                                              ���щ��                                                               ��BXYYYYZ                                                               �XXXYZZZZ                                                             YBXYZZZYYYY                                                           XBBYYYYZZ[ZYBXX                                                     �XAAAAAAABBXBBAB�                                                � XBAAAAAAAAAAAAAAA                                              �������BAAAAAA@AAAAAAAAA�                                              Ѡ�щ���AAAAAA��@AAAAA@��                                              蠈����AAAA���@��                                               �����щAAAA�������@��                                                  �ЉAAAA����������                                                    �Ј�AAAAA�����������                                                     �AAAAA������������                                                        �AAAAA������������                                                         �AAAA@������������                                                        �AAAA@�����������                                                         �AAA@�����������                                                         �AAA@������������                                                         �BAAA�����������                                                      XBA@�����������                                                    AA���������������                                              �AA���������������                                       Ј�AA�������������������                                     �����������뉈�������                                    ��������� ҉��������������                                    Ј���      �ss*++++++*++�                                   ���          s*++++++++++�                                                 ��r*++++++++++�                                                       �*��s*+++++++++++*�                                                     �++++��++++++++++++*�                                                    �+++��ь+++++++++++++�                                                  �++B�҉++++++++++***�                                                 ��+A�ӌ+++++++++***                                                �+++���++++++++*sss                                               �+++��s+++++++*�srs�sr                                             ��++++��s+++++*�ss���ssss�                                            �+++��s++++*sss������s����                                           ьB+++��r*+**�s����rrssssss�                                          BBBA��r***�s�   �srsss�ss�                                          A�������    ԋssssss��                                         �����       ԋssssss��                                        �������������         ыssssss�                                       �������������           ��������                                       �����������             �������                                       ���������                 ������                                       ꡣ�����                   �������                                        銣�                   ���                                       늣AA�                    鈊�                                        ���AA�                   ���A                                        ы�AA�                    ѡ�ABX                                       ���AA�                    �AAX                                       Ҋ��A��                    �AAA                                       �������                    �AAA�                                       ꊣ���                   �                                        ����                    ��A                                       늣�                     �A                                        ъ���                      �A�                                       ������                       ��                                        ꢤ��                        ���                                        ��                        �                                         颤�                        ��                                        ���                        �                                        ��                        ҡ�                                        ��                         �                                        Ң�                        Ѣ�                                       ꢤ�                      颤�                                      ����                   �                                      ����                   �艡���                                     ����                                                             �����                                                                 �                                                                 ��                                                                                                                         