��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       �                                                            �                                                            袣�                                                           ���                                                     �����                                                     �������                                                     ꡡ��� 눉���                                                      Ј��� �����                                                       뉠�����                                                   ꠠ��XBBAAA��                                                 ���XBBBBBBBBA���                                               ��XBBBBBBBXBBA���                                              ��AXBAAABBBYXBAA�                                       燈�       ТABAAAAAAABXXBAAAA�                                       ���      �AAAAAAAAAABBBBAAAA�                                       ����     ФAABBAA@AAABBAAAAAA�                                       ����   �AAAAAA��AAAAAAAAAAA�                                        袤  �AAAAAA����@AAAAAAAAAA�                                          ъ�ѢAAAAA����@@AAAAAAA�                                           Ң�AAAAA�����@@AAAA�                                           ���AAAAAAA������@A@��                                            �����AAAAA������@@@@��                                             Ҋ���AAAA��҈�������                                              ꋤ@A����҉��������                                               ҡ������҉���������                                                 щ�����ш��������������                                                      ��҉�������������                                                         ��҉������������                                                          ъ���������������                                                           Ѡ��������������                                                          ���������������                                                           ���������������                                                            Ҥ�������������                                                            ң�@�                                                           다@AAAAAAAA�                                                           ����@@AAAA@@��                                                          s***++AAAAAA����                                                         s**++++++++++++�                                                         r*�r++++++++++++�                                                       s**��s*++++++++++++�                                                      t++��s*++++++++++++�                                                     t++���*+++++++++++++�                                                    ��++���+++++++++++++++s                                                   s**�Ӊ++++++++++**+++*s                                                   r**��s++++*********�                                                 �*��s+++**�������                                                 �*���****�ssss����ssss�                                                �*���****ss�������rssss�                                               s��***ss������s�r                                               ���ss���   ��rsss                                              ��������     �rssss                                             ѣ������      �rsssss                                            �������s��        ��ssss�                                            ���������s�          ��sss��                                           ����������             ��ԉ���                                          ���������              ���늡�                                          ꣤������                ���뉡�                                          다���                   ��뉢�                                         ��AA                  ���X                                        ЊAABA                  ꊣAXY                                        ��ABB                   ��ABXY                                       �ABBB                   �AABYY                                      ��ABY�                    �ABBYY�                                     ��ABBA�                     �ABBY�                                      ѡ�ABA�                      ѣAABB�                                     ���AA�                      �AAB                                      ꢤAA                      ꡤAAB                                     ��AA                       �AB                                     ��AA                        �AB�                                     ��A�                          �A                                     ��A�                          �B                                     ѣ�A�                          ��                                     ��                           ��                                     �                            ���                                    ��                            ��                                    ��                           ���                                    �A                          ����                                  ��                         �������                                 衣�                     蠢�����뉉�                               뢣����                                                        ��������                                                            ����������                                                             ������                                                                                                                            