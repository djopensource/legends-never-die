��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                             ���                                                  ���                                                �����                                               Ј�����                                               鈉���                                               �뉊����    �                                             �ꉉ�����XY���������������                                   �ꈉ���BXYYZY���ꈈ���҈�������ABXZ                                   �鈉��AAAXX���������ꉊ������AABZ                                    �ꈊ��AA���������҈�������AAABYZ                                       鈉���A���������ꉉ������AAAAABY                                         ꉉ���������ꉉ������AAAAAA                                             ���������鈈������@AAAA                                                 룣��������뉉�����@A                                                ���������艉�������                                                 颤����ш�����������                                                  �����щ����щ����                                                  ѣ��������Ҥ�                                                   �����Ј����Т                                                  ����������Њ��                                                   �������Ј���������                                                   ���������������                                                    ъ��������������A                                                    �������������������                                                    ����ӈ�����������������                                                    ѣ����������������������                                                     ���������������������                                                     Ѥ������������Ӊ������                                                      ��������������ш�ꊡ�                                                       У������������ш�                                                        ��������������҉                                                            ��������������҉�                                                           ��������������ш�                                                          ���������������ъ�                                                          ꣣������������ҋ�                                                         Ћ������������rs*�                                                         Ӌ�����������*�                                                         �*������s**�                                                        �******�                                                        �**+++++*�                                                         �*++++++++*r�                                                         s*++++++++++r�                                                          �*++++++++*���                                                          �++++++++**�ѻ�                                                           �+++++++*�л�                                                           �+++++++*�҉                                                            �B++++++*���                                                            YAA+++*����                                                             �AAAA**�к��                                                            AAAAA��Ҋsr                                                            AAAAA����Ԋs�r                                                           AAA������sr�r                                                           XAA�������rrԻ�                                                          YA�����rss���                                                         ��������s���                                                         �����������҈                                                          �������   �����҈�                                                          ������    Ҋ��҈��                                                          鋢����   ���ꉉ�                                                         ����    ��ꈉ��                                                      ��   �ꈉ��AABY                                                    ��   ��ꉉ�AAAB                                                  ��    ���ꉉ����A�                                                ��    ������ꉉ����A�                                               ��      ���뉉���A�                                             ����             ��ꉊ���                                          �����                ��ꉊ���                                        ������                   �ꉊ��                                      �����                     ꉡ�                                     ����                        ꊣ�                                     ����                          ����                                     ����                         ����                                      ����                         ����                                       ����                        ����                                         ����                       ���                                          ѡ���                       ���                                          �����                       ���                                          ����                                                                    ����                                                                     �����                                                                    �����                                                                   �������                                                                 �����                                                                ����                                                               �                                                                                                             