��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                                                            щ���                                                             щ����                                                              ���鉡���                                                            ��҈�����                                                             ��ꈉ����                                                             ��뉉ꈉ����                                                              �����ш���                                                             ��������                                                           XAA���                                                          �YXXYYXAA�                                                             �YYYZZZYXAA�                                                           �YYYYZZZYYXBAX�                                                          XXYYZZYYXBAAAX                                                         �AAABBBBAAAAAAAAB                                                        �AAAAAAAA@@AAAAAB ��                                                �AAAAAAA@@@@@AAAA����                                                �AA@AAA��@@@AAA����                                                ��@@����@AAAAAA�����                                                �@@�������@AAAA@�����                                                ��������@AAAA@��렠���                                                 Ҥ��������AAAAAAA�����                                                    Т��������AAAAAA���                                                      ���������AAAAAA��                                                       룤������AAAAAA��                                                          ъ�������AAAAA�                                                           ���������@AAAA��                                                           ���������@AAAA�                                                          Ҋ�������@��AA                                                         щ����������@AA�                                                       ���������������AA                                                     �����������������AB                                             Ҥ����������������A����                                       �AA����������ꉉ������                                       Ҍ���@@���������ꉊ�����                                     �++**���������       ���                                     ��++++++++*��         Ј����                                     �++++++++++*****s                                              �++++++++++*�*+s                                                      �++++++++++r�+*�                                                      �+++++++++*�Ԍ++++��                                                      �+**++++++**sҊ+++++�                                                    �*+++++**r�ӌ+++++�                                                   ��*******t�щ�+++++�                                                 �sss***++*s�ы*+++�                                                ��sssrrs******��Ԍ*++��                                              �srrsrrrs�*****s�ҋ*++++�                                             �ssssr�rss�**��++++�                                            sssrrӺ��sssr�Ԍ++BA�                                           ssss�  ��sts�ҌAAAA                                          ssss�    �ss���AAA                                         sss��      ��st���                                        �ssss���        ��ss��������                                       �����s��          �ԉ�������                                      ��������               ҉�����                                      �������                 ꉉ����                                      �������                    ꣤���                                      щ�����                     ����                                     ������                     �A��                                    �BA����                     �AA���                                    XXAA��                      �AA��                                   YYBAA�                      AA���                                  �YBBA�                       �AA���                                  XBBBA�                        �A��                                  �ABBA�                         ���                                 �AAAAA��                          ����                                 �A��                           ����                                 �AA���                           ���                                 �AA��                             ���                                �AA��                              ����                                 �AA��                               ����                                �AA�                                ���                                ���                                ���                                ���                                ���                               ���                                 ���                               ���                                  �A��                              ����                               �AA�                             ����                            AA�                            ��������                            ����                           �����                                ��                          ��                                  �A                                                              �                                                              �렢��                                                                   ��         