��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ��                                                      YY                                                    YYYZZ                                                  YYZ[                                                 �YYZ[Z                                                �XYZZ[[                                               �ABYYZZ                                               �ꊣAABYY                                               ����ꉉ���AABYZ                                                 ������ꈉ����AABYZ�                                                 �����������҉�AABBYZZ�                                               �������������ӊAABBYZZZ�                                             �������������щ�AAABBXYYX                                            Ј�����������ш�AAAAAABB                                            �興�����������AAAAAAAA�                                           �����������������AAA@@AA�                                           ����������������҉AA@@�@���                                           ���ҊAA��������                                          ��            ѡ@���������                                                       �����������                                                      ���������뉢                                                     ����������뉋�                                                  ���������뉊��                                        Ј��        ��������뉉���                                       ����     �������ꈉ���A�                                      ����    ��������ꈉ���A��                                         Ј����  ��������҈�����A+�                                           ��������Ң�������҈����*+�                                           ��艡�������������ꈉ�*��                                             �ꊋ�����������������                                                щ������������rsss**�s�                                                 ш���������rrs***��ss                                                  ҈��������s*****��s�                                                     �ꈉ����++++++*�rs                                                       �҈��++++++*��s�                                                          ъ++++++*��s�                                                            �*+++++*���sr                                                           ��*++++*���ss                                                           ь***���ss�                                                           �***���ss�                                                           ����ss�                                                          �����ssr�                                                          ��������ssr��                                                          �A������ssrrӺ                                                         �A������ssr���                                                         ��������������                                                        �����눉�����                                                         ��������҈����                                                         ꣣����� �ꈈ���                                                         ������  ��ꉉ��                                                          ������   ��ꉊ�                                                         щ����  �҈����                                                       �����  �҈���                                                      ������  �҈��ABX�                                                     ������   ҈���ABXX                                                   ������   �ш���AAA�                                                  ������     �艢���                                                ������         ꉊ��                                               ������           �늣                                               ������             ҉���                                              ꡡ��               늢�                                            ꡡ��                 艡���                                          ꡊ��                    롤�                                         ꡡ��                     �                                        롡��                      ъ�                                        롊��                       뢤���                                        롊�                       뢣��                                         롊�                       ����                                         ����                       ��                                          ����                       ���                                           뢢��                      ��                                         ꢢ����                     鉉�                                       �������                    艈�                                     ��������                                                         ���������                                                             �����������                                                         �����������                                            