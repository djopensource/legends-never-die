��   �`]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ��                                                    YY                                                   ZZYYY                                                  [ZYY                                                Z[ZYY�                                               [[ZZYX�                                              ZZYYBA��                                             YYBAA����                                             ZYBAA����������                                             �ZYBAA�������������                                                �ZZYBBAA��������������                                                �ZZZYBBAA���������������                                              XYYXBBAAA����������������                                             BBAAAAAA�����������艉��                                            �AAAAAAAA�����������ꈈ��                                            �AA@@AAA������������������                                           ���@�@@AA������������������                                          ��������AA�����                                          ���������@��            ��                                          �����������                                                       ��뉊�������                                                      ꋉ�뉊�������                                                    ����눉�������                                                �����뉊������        Ј��                                      �A�����ꉊ�����     Ј��                                      ԌA�����ꉊ������    렠�                                     �+A������҈�������  �����                                        �+*������ꉊ������銣�����                                           ��*���ꈉ����������������                                           ���������������������                                             �s�**sssr��������������                                                ssҌ***srr�����������                                                  �sҌ*****s����������                                                   sr�*++++++��������                                                      �sӊ*++++++�����                                                        �sӉ*++++++��                                                           rs�Ԍ*+++++*�                                                              ss�ӌ*++++*��                                                             �ss�ӌ***��                                                             �ss�ы***�                                                            �ss�Њ�                                                            �rss�щ��                                                           ��rss��ԋ����                                                          ��rrss��ԋ��A�                                                          ���rssԉ����A�                                                         ����ԉ��������                                                          ��҈���눊���                                                         �ꈉ���҉�����                                                         ҉����� ꊢ�����                                                          щ�����  Ҋ����                                                        ������   Њ����                                                      �������  ������                                                      ������  �����                                                     �XBA�����  ꣤���                                                   XXBA�����   ������                                                  �AAA������   ������                                                ������     ������                                               �����         ������                                              ����           뢢���                                             �����             Ҋ����                                            ����               �����                                          ������                 �����                                         ����                    늊��                                        ��                     銡��                                        ���                      ъ���                                        ������                       Њ���                                         뢣��                       ����                                          롢�                       ����                                           ��                       ����                                           щ�                       ����                                           ��                      �����                                           艉�                     ъ�����                                          鈉�                    ъ�����                                                              ꡊ�����                                                               롊������                                                             銊��������                                                            �����������            